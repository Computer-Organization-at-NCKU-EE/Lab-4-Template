module Reg_M (
    input clk,
    input rst,
    input [31:0] alu_out_in,
    input [31:0] rs2_data_in, 
    input bubble_in,    
    output reg [31:0] alu_out_out,
    output reg [31:0] rs2_data_out,
    output reg bubble_out
);
    // TODO: finish Reg_M (memory stage) design
endmodule
